//1.Definicion del modulo y su I/O
//Dentro del parentesis se define el I/O

module _and (input a , input b , output c);
//2.Definicion de cables o componentes 
//3.Asignaciones , Instancias y conexiones 

assign c = a & b;

endmodule

